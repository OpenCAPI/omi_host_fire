-- $Id: tb_ln_dly1to4.vhdl 2455 2016-02-01 19:13:39Z lonny $
-- $URL: file:///afs/awd/projects/eclipz/c14/libs/fbc/.svnDB/p9ndd1/main/vhdl/tb_ln_dly1to4.vhdl $
-- @!Created with MAKESCH v.1.53
-- *!********************************************************************
-- *! (C) Copyright International Business Machines Corporation 2007-2013
-- *!           All Rights Reserved -- Property of IBM
-- *!                    *** IBM Confidential ***
-- *!********************************************************************
-- *! FILE NAME   :  tb_ln_dly1to4.vhdl
-- *! TITLE       :
-- *! DESCRIPTION : OpenCapi DL logic
-- *!
-- *!
-- *! OWNER NAME  :  Lambrecht, Lonny      (uid: lonny)
-- *! BACKUP NAME :  Ganfield, Paul        (uid: pag)
-- *!
-- *!********************************************************************
-- Revision History:
-- ----------------------------------------------------------------------
-- Version:|Author: | Date:  | Comment:
-- --------|--------|--------|-------------------------------------------
--         |lonny   |02/16/16| initial entry
-------------------------------------------------------------------------

---- MR_PARAMS -dec a -ri _din -clk opt_gckn -vd vdn -scan_ios -nolcbcntl -parse_subs
-- MR_PARAMS -dec a -ri _din -clk opt_gckn -vd vdn -parse_subs -sde tc_pbiooa_scan_diag_dc

-- Global VHDL language/common libraries:
library ibm, ieee, support, work;
 use ibm.std_ulogic_function_support.all;
 use ibm.std_ulogic_support.all;
 use ibm.synthesis_support.all;
 use ieee.std_logic_1164.all;
 use support.logic_support_pkg.all;

use ibm.std_ulogic_unsigned.all;

-- MAKE SCHEMATIC DIRECTIVES
-- MS_U



-- MAKEREGS IO DECLARATIONS START
Entity tb_ln_dly1to4 is port (

  delay                          : in  std_ulogic_vector(0 to 7);
  clock_in                       : in  std_ulogic;
  clk_in_phase                   : in  std_ulogic;
  lane_in_header                 : in  std_ulogic_vector(0 to 1);
  lane_in_data                   : in  std_ulogic_vector(0 to 63);
  lane_in_seq                    : in  std_ulogic_vector(0 to 5);
  lane_out                       : out std_ulogic_vector(0 to 15);


  inject_crc                     : in  std_ulogic;


---------------------------
-- clock controls
---------------------------

  opt_gckn                       : in  std_ulogic

);
 Attribute BLOCK_TYPE of tb_ln_dly1to4 : entity is leaf;
 Attribute BTR_NAME of tb_ln_dly1to4 : entity is "TB_LN_DLY1TO4";
 Attribute RECURSIVE_SYNTHESIS of tb_ln_dly1to4 : entity is 2;
 attribute pin_data of opt_gckn   : signal is "PIN_FUNCTION=/G_CLK/";


end tb_ln_dly1to4 ;
-- MAKEREGS IO DECLARATIONS END
-- MAKEREGS IO DECLARATIONS END
----------
Architecture tb_ln_dly1to4 of tb_ln_dly1to4 is


-- MAKEREGS SIGNAL DECLARATIONS START
-----------------------------------------------------------
-- Input and output signal declarations (including       --
-- scan signals) auto-generated by MAKEREGS version 309 --
-----------------------------------------------------------

-- Register signal declarations
  SIGNAL carryover_din, carryover_q : std_ulogic_vector(0 to 255);
  SIGNAL clk_cnt_din, clk_cnt_q : std_ulogic_vector(0 to 1);
  SIGNAL clock_din, clock_q : std_ulogic;
  SIGNAL delay_din, delay_q : std_ulogic_vector(0 to 7);
  SIGNAL init_din, init_q : std_ulogic;
  SIGNAL lane_in_din, lane_in_q : std_ulogic_vector(0 to 63);
  SIGNAL lane_out_din, lane_out_q : std_ulogic_vector(0 to 15);
  SIGNAL lfsr_din, lfsr_q : std_ulogic_vector(0 to 15);

-- Internal signal declarations
  SIGNAL act : std_ulogic;
  SIGNAL zeros : std_ulogic_vector(0 to 255);
  SIGNAL updated_lfsr : std_ulogic_vector(0 to 15);
  SIGNAL prev_in_data : std_ulogic_vector(0 to 63);
  SIGNAL prev_in_header : std_ulogic_vector(0 to 1);
  SIGNAL prev_in_seq : std_ulogic_vector(0 to 5);
  SIGNAL prev2_in_data : std_ulogic_vector(0 to 63);
  SIGNAL toggle : std_ulogic;
  SIGNAL seq_id : std_ulogic_vector(0 to 6);
  SIGNAL lane_in_int : std_ulogic_vector(0 to 15);

--  Enhancement to VS to help detect unused latch input/outputs
-- %VS_PORT_MAP c_nlat_scan.q out
-- %VS_PORT_MAP c_nlat_scan.qL1 out
-- %VS_PORT_MAP c_nlat_scan.data in
-- %VS_PORT_MAP c_nlat_scan.q out
-- %VS_PORT_MAP c_nlat_scan.qL1 out
-- %VS_PORT_MAP c_nlat_scan.data in
---------------------------------------------------------------
-- End auto-generated register and scan signal declarations  --
---------------------------------------------------------------
-- MAKEREGS SIGNAL DECLARATIONS END
attribute ANALYSIS_NOT_REFERENCED of carryover_q                           : signal is "<128:255>TRUE";
BEGIN
act                                          <= '1';
zeros (0 to 255)                             <= (others => '0');

init_din                     <= '1';
delay_din(0 to 7)            <= delay(0 to 7) when init_q = '0' else delay_q(0 to 7);
lfsr_din(0 to 15)            <= "1111111111111111"    when init_q = '0' else
                                updated_lfsr(0 to 15);

updated_lfsr(0)              <= lfsr_q(15);
updated_lfsr(1)              <= lfsr_q(0);
updated_lfsr(2)              <= lfsr_q(1) xor lfsr_q(15);  -- 
updated_lfsr(3)              <= lfsr_q(2) xor lfsr_q(15);
updated_lfsr(4)              <= lfsr_q(3);
updated_lfsr(5)              <= lfsr_q(4) xor lfsr_q(15);
updated_lfsr(6 to 15)        <= lfsr_q(5 to 14);

clock_din                    <= clock_in;

-- MAKESCH GENERATED
    prev : entity work.tb_ln_dly1to4_4x
    port map (
        lane_in_data (0 to 63)         => lane_in_data (0 to 63)         , -- OVR: tb_ln_dly1to4_4x(prev)
        lane_in_header (0 to 1)        => lane_in_header (0 to 1)        , -- OVR: tb_ln_dly1to4_4x(prev)
        lane_in_seq (0 to 5)           => lane_in_seq (0 to 5)           , -- OVR: tb_ln_dly1to4_4x(prev)
        prev_in_data (0 to 63)         => prev_in_data (0 to 63)         , -- OVD: tb_ln_dly1to4_4x(prev)
        prev_in_header (0 to 1)        => prev_in_header (0 to 1)        , -- OVD: tb_ln_dly1to4_4x(prev)
        prev_in_seq (0 to 5)           => prev_in_seq (0 to 5)           , -- OVD: tb_ln_dly1to4_4x(prev)
        prev2_in_data (0 to 63)        => prev2_in_data (0 to 63)        , -- OVD: tb_ln_dly1to4_4x(prev)
        opt_gckn                       => clock_in                         -- OVR: tb_ln_dly1to4_4x(prev)
    ) ;
-- MAKESCH GENERATED ENDS

toggle                       <= prev_in_seq(0 to 5) = lane_in_seq(0 to 5);
seq_id(0 to 6)             <= lane_in_seq(0 to 5) & toggle;

with seq_id(0 to 6) select
lane_in_din(0 to 63)         <=                           lane_in_header(0 to 1) & lane_in_data(0 to 61)  when "0000000",
                                prev_in_data(62 to 63)  & lane_in_header(0 to 1) & lane_in_data(0 to 59)  when "0000001",
                                prev_in_data(60 to 63)  & lane_in_header(0 to 1) & lane_in_data(0 to 57)  when "0000010",
                                prev_in_data(58 to 63)  & lane_in_header(0 to 1) & lane_in_data(0 to 55)  when "0000011",
                                prev_in_data(56 to 63)  & lane_in_header(0 to 1) & lane_in_data(0 to 53)  when "0000100",
                                prev_in_data(54 to 63)  & lane_in_header(0 to 1) & lane_in_data(0 to 51)  when "0000101",
                                prev_in_data(52 to 63)  & lane_in_header(0 to 1) & lane_in_data(0 to 49)  when "0000110",
                                prev_in_data(50 to 63)  & lane_in_header(0 to 1) & lane_in_data(0 to 47)  when "0000111",
                                prev_in_data(48 to 63)  & lane_in_header(0 to 1) & lane_in_data(0 to 45)  when "0001000",
                                prev_in_data(46 to 63)  & lane_in_header(0 to 1) & lane_in_data(0 to 43)  when "0001001",
                                prev_in_data(44 to 63)  & lane_in_header(0 to 1) & lane_in_data(0 to 41)  when "0001010",
                                prev_in_data(42 to 63)  & lane_in_header(0 to 1) & lane_in_data(0 to 39)  when "0001011",
                                prev_in_data(40 to 63)  & lane_in_header(0 to 1) & lane_in_data(0 to 37)  when "0001100",
                                prev_in_data(38 to 63)  & lane_in_header(0 to 1) & lane_in_data(0 to 35)  when "0001101",
                                prev_in_data(36 to 63)  & lane_in_header(0 to 1) & lane_in_data(0 to 33)  when "0001110",
                                prev_in_data(34 to 63)  & lane_in_header(0 to 1) & lane_in_data(0 to 31)  when "0001111",
                                prev_in_data(32 to 63)  & lane_in_header(0 to 1) & lane_in_data(0 to 29)  when "0010000",
                                prev_in_data(30 to 63)  & lane_in_header(0 to 1) & lane_in_data(0 to 27)  when "0010001",
                                prev_in_data(28 to 63)  & lane_in_header(0 to 1) & lane_in_data(0 to 25)  when "0010010",
                                prev_in_data(26 to 63)  & lane_in_header(0 to 1) & lane_in_data(0 to 23)  when "0010011",
                                prev_in_data(24 to 63)  & lane_in_header(0 to 1) & lane_in_data(0 to 21)  when "0010100",
                                prev_in_data(22 to 63)  & lane_in_header(0 to 1) & lane_in_data(0 to 19)  when "0010101",
                                prev_in_data(20 to 63)  & lane_in_header(0 to 1) & lane_in_data(0 to 17)  when "0010110",
                                prev_in_data(18 to 63)  & lane_in_header(0 to 1) & lane_in_data(0 to 15)  when "0010111",
                                prev_in_data(16 to 63)  & lane_in_header(0 to 1) & lane_in_data(0 to 13)  when "0011000",
                                prev_in_data(14 to 63)  & lane_in_header(0 to 1) & lane_in_data(0 to 11)  when "0011001",
                                prev_in_data(12 to 63)  & lane_in_header(0 to 1) & lane_in_data(0 to  9)  when "0011010",
                                prev_in_data(10 to 63)  & lane_in_header(0 to 1) & lane_in_data(0 to  7)  when "0011011",
                                prev_in_data( 8 to 63)  & lane_in_header(0 to 1) & lane_in_data(0 to  5)  when "0011100",
                                prev_in_data( 6 to 63)  & lane_in_header(0 to 1) & lane_in_data(0 to  3)  when "0011101",
                                prev_in_data( 4 to 63)  & lane_in_header(0 to 1) & lane_in_data(0 to  1)  when "0011110",
                                prev_in_data( 2 to 63)  & lane_in_header(0 to 1)                          when "0011111",
                                prev_in_data( 0 to 63)                                                    when "0100000",
                                                          prev_in_header(0 to 1) & prev_in_data(0 to 61)  when "0100001",
                                prev2_in_data(62 to 63) & prev_in_header(0 to 1) & prev_in_data(0 to 59)  when "0100010",
                                prev2_in_data(60 to 63) & prev_in_header(0 to 1) & prev_in_data(0 to 57)  when "0100011",
                                prev2_in_data(58 to 63) & prev_in_header(0 to 1) & prev_in_data(0 to 55)  when "0100100",
                                prev2_in_data(56 to 63) & prev_in_header(0 to 1) & prev_in_data(0 to 53)  when "0100101",
                                prev2_in_data(54 to 63) & prev_in_header(0 to 1) & prev_in_data(0 to 51)  when "0100110",
                                prev2_in_data(52 to 63) & prev_in_header(0 to 1) & prev_in_data(0 to 49)  when "0100111",
                                prev2_in_data(50 to 63) & prev_in_header(0 to 1) & prev_in_data(0 to 47)  when "0101000",
                                prev2_in_data(48 to 63) & prev_in_header(0 to 1) & prev_in_data(0 to 45)  when "0101001",
                                prev2_in_data(46 to 63) & prev_in_header(0 to 1) & prev_in_data(0 to 43)  when "0101010",
                                prev2_in_data(44 to 63) & prev_in_header(0 to 1) & prev_in_data(0 to 41)  when "0101011",
                                prev2_in_data(42 to 63) & prev_in_header(0 to 1) & prev_in_data(0 to 39)  when "0101100",
                                prev2_in_data(40 to 63) & prev_in_header(0 to 1) & prev_in_data(0 to 37)  when "0101101",
                                prev2_in_data(38 to 63) & prev_in_header(0 to 1) & prev_in_data(0 to 35)  when "0101110",
                                prev2_in_data(36 to 63) & prev_in_header(0 to 1) & prev_in_data(0 to 33)  when "0101111",
                                prev2_in_data(34 to 63) & prev_in_header(0 to 1) & prev_in_data(0 to 31)  when "0110000",
                                prev2_in_data(32 to 63) & prev_in_header(0 to 1) & prev_in_data(0 to 29)  when "0110001",
                                prev2_in_data(30 to 63) & prev_in_header(0 to 1) & prev_in_data(0 to 27)  when "0110010",
                                prev2_in_data(28 to 63) & prev_in_header(0 to 1) & prev_in_data(0 to 25)  when "0110011",
                                prev2_in_data(26 to 63) & prev_in_header(0 to 1) & prev_in_data(0 to 23)  when "0110100",
                                prev2_in_data(24 to 63) & prev_in_header(0 to 1) & prev_in_data(0 to 21)  when "0110101",
                                prev2_in_data(22 to 63) & prev_in_header(0 to 1) & prev_in_data(0 to 19)  when "0110110",
                                prev2_in_data(20 to 63) & prev_in_header(0 to 1) & prev_in_data(0 to 17)  when "0110111",
                                prev2_in_data(18 to 63) & prev_in_header(0 to 1) & prev_in_data(0 to 15)  when "0111000",
                                prev2_in_data(16 to 63) & prev_in_header(0 to 1) & prev_in_data(0 to 13)  when "0111001",
                                prev2_in_data(14 to 63) & prev_in_header(0 to 1) & prev_in_data(0 to 11)  when "0111010",
                                prev2_in_data(12 to 63) & prev_in_header(0 to 1) & prev_in_data(0 to  9)  when "0111011",
                                prev2_in_data(10 to 63) & prev_in_header(0 to 1) & prev_in_data(0 to  7)  when "0111100",
                                prev2_in_data( 8 to 63) & prev_in_header(0 to 1) & prev_in_data(0 to  5)  when "0111101",
                                prev2_in_data( 6 to 63) & prev_in_header(0 to 1) & prev_in_data(0 to  3)  when "0111110",
                                prev2_in_data( 4 to 63) & prev_in_header(0 to 1) & prev_in_data(0 to  1)  when "0111111",
                                prev2_in_data( 2 to 63) & prev_in_header(0 to 1)                          when "1000000",
                                prev2_in_data( 0 to 63)                                                   when others;
                                

lane_in_int(0 to 15)         <= lane_in_q( 0 to 15) when clk_cnt_q(0 to 1) = "00" else
                                lane_in_q(16 to 31) when clk_cnt_q(0 to 1) = "01" else
                                lane_in_q(32 to 47) when clk_cnt_q(0 to 1) = "10" else
                                lane_in_q(48 to 63);

clk_cnt_din(0 to 1)          <= "00" when (clock_in = '0' and clock_q = '1' and clk_in_phase = '0') else 
                                "11" when (clock_in = '0' and clock_q = '1' and clk_in_phase = '1') else 
                                clk_cnt_q(0 to 1) + 1;

--lane_out(0 to 15)                            <= lane_out_q(0 to 15);
lane_out(0 to 15)                            <= lane_out_q(0 to 15) when inject_crc = '0' else (lane_out_q(0 to 14) & not lane_out_q(15));

with delay_q(0 to 7) select
lane_out_din(0 to 15)                        <=                        lane_in_int(0 to 15)     when "00000000",
                                                carryover_q(0)       & lane_in_int(0 to 14)     when "00000001",
                                                carryover_q(0 to  1) & lane_in_int(0 to 13)     when "00000010",
                                                carryover_q(0 to  2) & lane_in_int(0 to 12)     when "00000011",
                                                carryover_q(0 to  3) & lane_in_int(0 to 11)     when "00000100",
                                                carryover_q(0 to  4) & lane_in_int(0 to 10)     when "00000101",
                                                carryover_q(0 to  5) & lane_in_int(0 to  9)     when "00000110",
                                                carryover_q(0 to  6) & lane_in_int(0 to  8)     when "00000111",
                                                carryover_q(0 to  7) & lane_in_int(0 to  7)     when "00001000",
                                                carryover_q(0 to  8) & lane_in_int(0 to  6)     when "00001001",
                                                carryover_q(0 to  9) & lane_in_int(0 to  5)     when "00001010",
                                                carryover_q(0 to 10) & lane_in_int(0 to  4)     when "00001011",
                                                carryover_q(0 to 11) & lane_in_int(0 to  3)     when "00001100",
                                                carryover_q(0 to 12) & lane_in_int(0 to  2)     when "00001101",
                                                carryover_q(0 to 13) & lane_in_int(0 to  1)     when "00001110",
                                                carryover_q(0 to 14) & lane_in_int(0)           when "00001111",
                                                zeros(0 to 15)                                  when "11111110",
                                                lfsr_q(0 to 15)                                 when "11111111",
                                                carryover_q(0 to 15)                            when others;

with delay_q(0 to 7) select
carryover_din(0 to 255)                      <=                                                  zeros(0 to 255)     when "00000000",
                                                                         lane_in_int(15)       & zeros(0 to 254)     when "00000001",
                                                                         lane_in_int(14 to 15) & zeros(0 to 253)     when "00000010",
                                                                         lane_in_int(13 to 15) & zeros(0 to 252)     when "00000011",
                                                                         lane_in_int(12 to 15) & zeros(0 to 251)     when "00000100",
                                                                         lane_in_int(11 to 15) & zeros(0 to 250)     when "00000101",
                                                                         lane_in_int(10 to 15) & zeros(0 to 249)     when "00000110",
                                                                         lane_in_int( 9 to 15) & zeros(0 to 248)     when "00000111",
                                                                         lane_in_int( 8 to 15) & zeros(0 to 247)     when "00001000",
                                                                         lane_in_int( 7 to 15) & zeros(0 to 246)     when "00001001",
                                                                         lane_in_int( 6 to 15) & zeros(0 to 245)     when "00001010",
                                                                         lane_in_int( 5 to 15) & zeros(0 to 244)     when "00001011",
                                                                         lane_in_int( 4 to 15) & zeros(0 to 243)     when "00001100",
                                                                         lane_in_int( 3 to 15) & zeros(0 to 242)     when "00001101",
                                                                         lane_in_int( 2 to 15) & zeros(0 to 241)     when "00001110",
                                                                         lane_in_int( 1 to 15) & zeros(0 to 240)     when "00001111",
                                                                         lane_in_int( 0 to 15) & zeros(0 to 239)     when "00010000",
                                                carryover_q(16)        & lane_in_int( 0 to 15) & zeros(0 to 238)     when "00010001",
                                                carryover_q(16 to  17) & lane_in_int( 0 to 15) & zeros(0 to 237)     when "00010010",
                                                carryover_q(16 to  18) & lane_in_int( 0 to 15) & zeros(0 to 236)     when "00010011",
                                                carryover_q(16 to  19) & lane_in_int( 0 to 15) & zeros(0 to 235)     when "00010100",
                                                carryover_q(16 to  20) & lane_in_int( 0 to 15) & zeros(0 to 234)     when "00010101",
                                                carryover_q(16 to  21) & lane_in_int( 0 to 15) & zeros(0 to 233)     when "00010110",
                                                carryover_q(16 to  22) & lane_in_int( 0 to 15) & zeros(0 to 232)     when "00010111",
                                                carryover_q(16 to  23) & lane_in_int( 0 to 15) & zeros(0 to 231)     when "00011000",
                                                carryover_q(16 to  24) & lane_in_int( 0 to 15) & zeros(0 to 230)     when "00011001",
                                                carryover_q(16 to  25) & lane_in_int( 0 to 15) & zeros(0 to 229)     when "00011010",
                                                carryover_q(16 to  26) & lane_in_int( 0 to 15) & zeros(0 to 228)     when "00011011",
                                                carryover_q(16 to  27) & lane_in_int( 0 to 15) & zeros(0 to 227)     when "00011100",
                                                carryover_q(16 to  28) & lane_in_int( 0 to 15) & zeros(0 to 226)     when "00011101",
                                                carryover_q(16 to  29) & lane_in_int( 0 to 15) & zeros(0 to 225)     when "00011110",
                                                carryover_q(16 to  30) & lane_in_int( 0 to 15) & zeros(0 to 224)     when "00011111",
                                                carryover_q(16 to  31) & lane_in_int( 0 to 15) & zeros(0 to 223)     when "00100000",
                                                carryover_q(16 to  32) & lane_in_int( 0 to 15) & zeros(0 to 222)     when "00100001",
                                                carryover_q(16 to  33) & lane_in_int( 0 to 15) & zeros(0 to 221)     when "00100010",
                                                carryover_q(16 to  34) & lane_in_int( 0 to 15) & zeros(0 to 220)     when "00100011",
                                                carryover_q(16 to  35) & lane_in_int( 0 to 15) & zeros(0 to 219)     when "00100100",
                                                carryover_q(16 to  36) & lane_in_int( 0 to 15) & zeros(0 to 218)     when "00100101",
                                                carryover_q(16 to  37) & lane_in_int( 0 to 15) & zeros(0 to 217)     when "00100110",
                                                carryover_q(16 to  38) & lane_in_int( 0 to 15) & zeros(0 to 216)     when "00100111",
                                                carryover_q(16 to  39) & lane_in_int( 0 to 15) & zeros(0 to 215)     when "00101000",
                                                carryover_q(16 to  40) & lane_in_int( 0 to 15) & zeros(0 to 214)     when "00101001",
                                                carryover_q(16 to  41) & lane_in_int( 0 to 15) & zeros(0 to 213)     when "00101010",
                                                carryover_q(16 to  42) & lane_in_int( 0 to 15) & zeros(0 to 212)     when "00101011",
                                                carryover_q(16 to  43) & lane_in_int( 0 to 15) & zeros(0 to 211)     when "00101100",
                                                carryover_q(16 to  44) & lane_in_int( 0 to 15) & zeros(0 to 210)     when "00101101",
                                                carryover_q(16 to  45) & lane_in_int( 0 to 15) & zeros(0 to 209)     when "00101110",
                                                carryover_q(16 to  46) & lane_in_int( 0 to 15) & zeros(0 to 208)     when "00101111",
                                                carryover_q(16 to  47) & lane_in_int( 0 to 15) & zeros(0 to 207)     when "00110000",
                                                carryover_q(16 to  48) & lane_in_int( 0 to 15) & zeros(0 to 206)     when "00110001",
                                                carryover_q(16 to  49) & lane_in_int( 0 to 15) & zeros(0 to 205)     when "00110010",
                                                carryover_q(16 to  50) & lane_in_int( 0 to 15) & zeros(0 to 204)     when "00110011",
                                                carryover_q(16 to  51) & lane_in_int( 0 to 15) & zeros(0 to 203)     when "00110100",
                                                carryover_q(16 to  52) & lane_in_int( 0 to 15) & zeros(0 to 202)     when "00110101",
                                                carryover_q(16 to  53) & lane_in_int( 0 to 15) & zeros(0 to 201)     when "00110110",
                                                carryover_q(16 to  54) & lane_in_int( 0 to 15) & zeros(0 to 200)     when "00110111",
                                                carryover_q(16 to  55) & lane_in_int( 0 to 15) & zeros(0 to 199)     when "00111000",
                                                carryover_q(16 to  56) & lane_in_int( 0 to 15) & zeros(0 to 198)     when "00111001",
                                                carryover_q(16 to  57) & lane_in_int( 0 to 15) & zeros(0 to 197)     when "00111010",
                                                carryover_q(16 to  58) & lane_in_int( 0 to 15) & zeros(0 to 196)     when "00111011",
                                                carryover_q(16 to  59) & lane_in_int( 0 to 15) & zeros(0 to 195)     when "00111100",
                                                carryover_q(16 to  60) & lane_in_int( 0 to 15) & zeros(0 to 194)     when "00111101",
                                                carryover_q(16 to  61) & lane_in_int( 0 to 15) & zeros(0 to 193)     when "00111110",
                                                carryover_q(16 to  62) & lane_in_int( 0 to 15) & zeros(0 to 192)     when "00111111",
                                                carryover_q(16 to  63) & lane_in_int( 0 to 15) & zeros(0 to 191)     when "01000000",
                                                carryover_q(16 to  64) & lane_in_int( 0 to 15) & zeros(0 to 190)     when "01000001",
                                                carryover_q(16 to  65) & lane_in_int( 0 to 15) & zeros(0 to 189)     when "01000010",
                                                carryover_q(16 to  66) & lane_in_int( 0 to 15) & zeros(0 to 188)     when "01000011",
                                                carryover_q(16 to  67) & lane_in_int( 0 to 15) & zeros(0 to 187)     when "01000100",
                                                carryover_q(16 to  68) & lane_in_int( 0 to 15) & zeros(0 to 186)     when "01000101",
                                                carryover_q(16 to  69) & lane_in_int( 0 to 15) & zeros(0 to 185)     when "01000110",
                                                carryover_q(16 to  70) & lane_in_int( 0 to 15) & zeros(0 to 184)     when "01000111",
                                                carryover_q(16 to  71) & lane_in_int( 0 to 15) & zeros(0 to 183)     when "01001000",
                                                carryover_q(16 to  72) & lane_in_int( 0 to 15) & zeros(0 to 182)     when "01001001",
                                                carryover_q(16 to  73) & lane_in_int( 0 to 15) & zeros(0 to 181)     when "01001010",
                                                carryover_q(16 to  74) & lane_in_int( 0 to 15) & zeros(0 to 180)     when "01001011",
                                                carryover_q(16 to  75) & lane_in_int( 0 to 15) & zeros(0 to 179)     when "01001100",
                                                carryover_q(16 to  76) & lane_in_int( 0 to 15) & zeros(0 to 178)     when "01001101",
                                                carryover_q(16 to  77) & lane_in_int( 0 to 15) & zeros(0 to 177)     when "01001110",
                                                carryover_q(16 to  78) & lane_in_int( 0 to 15) & zeros(0 to 176)     when "01001111",
                                                carryover_q(16 to  79) & lane_in_int( 0 to 15) & zeros(0 to 175)     when "01010000",
                                                carryover_q(16 to  80) & lane_in_int( 0 to 15) & zeros(0 to 174)     when "01010001",
                                                carryover_q(16 to  81) & lane_in_int( 0 to 15) & zeros(0 to 173)     when "01010010",
                                                carryover_q(16 to  82) & lane_in_int( 0 to 15) & zeros(0 to 172)     when "01010011",
                                                carryover_q(16 to  83) & lane_in_int( 0 to 15) & zeros(0 to 171)     when "01010100",
                                                carryover_q(16 to  84) & lane_in_int( 0 to 15) & zeros(0 to 170)     when "01010101",
                                                carryover_q(16 to  85) & lane_in_int( 0 to 15) & zeros(0 to 169)     when "01010110",
                                                carryover_q(16 to  86) & lane_in_int( 0 to 15) & zeros(0 to 168)     when "01010111",
                                                carryover_q(16 to  87) & lane_in_int( 0 to 15) & zeros(0 to 167)     when "01011000",
                                                carryover_q(16 to  88) & lane_in_int( 0 to 15) & zeros(0 to 166)     when "01011001",
                                                carryover_q(16 to  89) & lane_in_int( 0 to 15) & zeros(0 to 165)     when "01011010",
                                                carryover_q(16 to  90) & lane_in_int( 0 to 15) & zeros(0 to 164)     when "01011011",
                                                carryover_q(16 to  91) & lane_in_int( 0 to 15) & zeros(0 to 163)     when "01011100",
                                                carryover_q(16 to  92) & lane_in_int( 0 to 15) & zeros(0 to 162)     when "01011101",
                                                carryover_q(16 to  93) & lane_in_int( 0 to 15) & zeros(0 to 161)     when "01011110",
                                                carryover_q(16 to  94) & lane_in_int( 0 to 15) & zeros(0 to 160)     when "01011111",
                                                carryover_q(16 to  95) & lane_in_int( 0 to 15) & zeros(0 to 159)     when "01100000",
                                                carryover_q(16 to  96) & lane_in_int( 0 to 15) & zeros(0 to 158)     when "01100001",
                                                carryover_q(16 to  97) & lane_in_int( 0 to 15) & zeros(0 to 157)     when "01100010",
                                                carryover_q(16 to  98) & lane_in_int( 0 to 15) & zeros(0 to 156)     when "01100011",
                                                carryover_q(16 to  99) & lane_in_int( 0 to 15) & zeros(0 to 155)     when "01100100",
                                                carryover_q(16 to 100) & lane_in_int( 0 to 15) & zeros(0 to 154)     when "01100101",
                                                carryover_q(16 to 101) & lane_in_int( 0 to 15) & zeros(0 to 153)     when "01100110",
                                                carryover_q(16 to 102) & lane_in_int( 0 to 15) & zeros(0 to 152)     when "01100111",
                                                carryover_q(16 to 103) & lane_in_int( 0 to 15) & zeros(0 to 151)     when "01101000",
                                                carryover_q(16 to 104) & lane_in_int( 0 to 15) & zeros(0 to 150)     when "01101001",
                                                carryover_q(16 to 105) & lane_in_int( 0 to 15) & zeros(0 to 149)     when "01101010",
                                                carryover_q(16 to 106) & lane_in_int( 0 to 15) & zeros(0 to 148)     when "01101011",
                                                carryover_q(16 to 107) & lane_in_int( 0 to 15) & zeros(0 to 147)     when "01101100",
                                                carryover_q(16 to 108) & lane_in_int( 0 to 15) & zeros(0 to 146)     when "01101101",
                                                carryover_q(16 to 109) & lane_in_int( 0 to 15) & zeros(0 to 145)     when "01101110",
                                                carryover_q(16 to 110) & lane_in_int( 0 to 15) & zeros(0 to 144)     when "01101111",
                                                carryover_q(16 to 111) & lane_in_int( 0 to 15) & zeros(0 to 143)     when "01110000",
                                                carryover_q(16 to 112) & lane_in_int( 0 to 15) & zeros(0 to 142)     when "01110001",
                                                carryover_q(16 to 113) & lane_in_int( 0 to 15) & zeros(0 to 141)     when "01110010",
                                                carryover_q(16 to 114) & lane_in_int( 0 to 15) & zeros(0 to 140)     when "01110011",
                                                carryover_q(16 to 115) & lane_in_int( 0 to 15) & zeros(0 to 139)     when "01110100",
                                                carryover_q(16 to 116) & lane_in_int( 0 to 15) & zeros(0 to 138)     when "01110101",
                                                carryover_q(16 to 117) & lane_in_int( 0 to 15) & zeros(0 to 137)     when "01110110",
                                                carryover_q(16 to 118) & lane_in_int( 0 to 15) & zeros(0 to 136)     when "01110111",
                                                carryover_q(16 to 119) & lane_in_int( 0 to 15) & zeros(0 to 135)     when "01111000",
                                                carryover_q(16 to 120) & lane_in_int( 0 to 15) & zeros(0 to 134)     when "01111001",
                                                carryover_q(16 to 121) & lane_in_int( 0 to 15) & zeros(0 to 133)     when "01111010",
                                                carryover_q(16 to 122) & lane_in_int( 0 to 15) & zeros(0 to 132)     when "01111011",
                                                carryover_q(16 to 123) & lane_in_int( 0 to 15) & zeros(0 to 131)     when "01111100",
                                                carryover_q(16 to 124) & lane_in_int( 0 to 15) & zeros(0 to 130)     when "01111101",
                                                carryover_q(16 to 125) & lane_in_int( 0 to 15) & zeros(0 to 129)     when "01111110",
                                                carryover_q(16 to 126) & lane_in_int( 0 to 15) & zeros(0 to 128)     when "01111111",
                                                carryover_q(16 to 127) & lane_in_int( 0 to 15) & zeros(0 to 127)     when others;

  carryoverq: entity work.fire_morph_dff
    generic map (width => 256)
    port map(gckn            => opt_gckn,
             e               => act,
             d               => carryover_din(0 to 255),
             q               => carryover_q(0 to 255));

  clk_cntq: entity work.fire_morph_dff
    generic map (width => 2)
    port map(gckn            => opt_gckn,
             e               => act,
             d               => clk_cnt_din(0 to 1),
             q               => clk_cnt_q(0 to 1));

  clockq: entity work.fire_morph_dff
    generic map (width => 1)
    port map(gckn            => opt_gckn,
             e               => act,
             d(0)            => clock_din,
             q(0)            => clock_q );

  delayq: entity work.fire_morph_dff
    generic map (width => 8)
    port map(gckn            => opt_gckn,
             e               => act,
             d               => delay_din(0 to 7),
             q               => delay_q(0 to 7));

  initq: entity work.fire_morph_dff
    generic map (width => 1)
    port map(gckn            => opt_gckn,
             e               => act,
             d(0)            => init_din,
             q(0)            => init_q );

  lane_inq: entity work.fire_morph_dff
    generic map (width => 64)
    port map(gckn            => opt_gckn,
             e               => act,
             d               => lane_in_din(0 to 63),
             q               => lane_in_q(0 to 63));

  lane_outq: entity work.fire_morph_dff
    generic map (width => 16)
    port map(gckn            => opt_gckn,
             e               => act,
             d               => lane_out_din(0 to 15),
             q               => lane_out_q(0 to 15));

  lfsrq: entity work.fire_morph_dff
    generic map (width => 16)
    port map(gckn            => opt_gckn,
             e               => act,
             d               => lfsr_din(0 to 15),
             q               => lfsr_q(0 to 15));
End tb_ln_dly1to4;
